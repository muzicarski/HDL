`ifndef FIFO_TYPES_PKG_SV
 `define FIFO_TYPES_PKG_SV


typedef enum {READ = 0, WRITE = 1, RW = 2} op_t;




`endif
